-------------------------------------------------------------------------
-- Engineer    : Golovachenko Victor
--
-- Create Date : 13.01.2016 17:12:50
-- Module Name : ust_def
--
-- Description :
--
-------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

package ust_def is

constant C_PKT_TYPE_VIDEO : natural := 1;

constant C_VIDEO_PKT_HEADER_BYTECOUNT : natural := 16;

end package ust_def;

